-- Sol Ayelen Cataldo 
-- Voltimetro que es la suma de todos los caracteres
entity voltimetro_tb is
end entity voltimetro_tb;

architecture voltimetro_tb_arq of voltimetro_tb is

begin
	
end architecture voltimetro_tb_arq;
